module rom(
	input [15:0] Adds,
	output wire [31:0] Inst
);
//escrever programa aqui em linguagem de máquina
endmodule